typedef uvm_sequencer#(unpacker_transaction) unpacker_sequencer;
