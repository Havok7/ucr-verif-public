typedef uvm_sequencer#(c3po_transaction) c3po_sequencer;
